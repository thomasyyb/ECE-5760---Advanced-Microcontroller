module solver (

);

endmodule 

