module compute_harmonic (
    input logic n,
    input logic L,
    input logic K,
);




endmodule 